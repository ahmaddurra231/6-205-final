//this module is currently not being used 
module address_generator #(parameter ADDR_WIDTH = 8)(
  input wire clk_in,
  input wire rst_in,
  output logic [7:0] address_out
);
  
endmodule